<!doctype html>
	<html lang="sv">
		<head>
			<meta charset="utf-8" />
			<title>409 Conflict</title>
			<style type="text/css">
				html {
					height: 100%;
				}
				body {
					color: #3A3A3A;
					font-family: Arial, sans-serif;
					font-size: 1.2em;
					background-color: #F6F6F6;
					padding: 0px;
					margin: 0px;
					height: 100%;
					overflow: hidden;
				}
				h1 {
					font-family: Arial, sans-serif;	
					font-weight: 900;
					font-size: 3em;
					color: #002e54;
					text-align: center;
				}
				h2 {
					font-family: Arial, sans-serif;	
					font-weight: bold;
					font-size: 1em;
					color: #777;
					text-align: left;	
				}
				h3 {
					font-family: Arial, sans-serif;	
					font-weight: bold;
					font-size: 1em;
					color: #777;
					text-align: left;		
				}
				a {
					color: #002e54;
					text-decoration: none;
				}
				a:hover {
					color: #006DB2;
				}
				#wrapper {
					width: 100%;
					height: 100%;
				}
				#content {
					width: 600px;
					height: 100%;
					padding: 40px 20px;
					margin: auto;
					background-color: #fff;
					border-left: 1px solid #cccccc;
					border-right: 1px solid #cccccc;
				}
				img#wikialogo {
					width: 50%;
					margin: 0px auto;
					display: block;
				}
				div.links {
					margin-top: 30px;
					font-size: 0.8em;
				}
				div.technical {
					margin-top: 60px;
					font-size: 0.6em;
					color: #777;
				}

			</style>
			<!--[if IE]>
			<script src="http://html5shiv.googlecode.com/svn/trunk/html5.js"></script>
			<![endif]-->
		</head>
		<body>
			<div id="wrapper">
				<div id="content">
					<img src="http://upload.wikimedia.org/wikipedia/commons/1/17/Wikia_Logo.svg" id="wikialogo"/>
					<div class="friendly">
						<h1>We are sorry!</h1>
						<p>There is some kind of conflict. Please check the URL for mistakes.</p>
					</div>
					<div class="links">
						For more info and updates check out our <a href="https://twitter.com/Wikia">Twitter Feed</a>.
					</div>
					<div class="technical">
						<h2>Technical explanation for geeks and administrators:</h2>
						<h3>409 Conflict</h3>
						<p>The request could not be completed due to a conflict with the current state of the resource. This code is only allowed in situations where it is expected that the user might be able to resolve the conflict and resubmit the request.</p>
					</div>
			</div> <!-- #content -->
		</div> <!-- #wrapper -->
	</body>
</html>