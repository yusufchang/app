<!doctype html>
	<html lang="sv">
		<head>
			<meta charset="utf-8" />
			<title>502 Bad Gateaway</title>
			<style type="text/css">
				html {
					height: 100%;
				}
				body {
					color: #3A3A3A;
					font-family: Arial, sans-serif;
					font-size: 1.2em;
					background-color: #F6F6F6;
					padding: 0px;
					margin: 0px;
					height: 100%;
					overflow: hidden;
				}
				h1 {
					font-family: Arial, sans-serif;	
					font-weight: 900;
					font-size: 3em;
					color: #002e54;
					text-align: center;
				}
				h2 {
					font-family: Arial, sans-serif;	
					font-weight: bold;
					font-size: 1em;
					color: #777;
					text-align: left;	
				}
				h3 {
					font-family: Arial, sans-serif;	
					font-weight: bold;
					font-size: 1em;
					color: #777;
					text-align: left;		
				}
				a {
					color: #002e54;
					text-decoration: none;
				}
				a:hover {
					color: #006DB2;
				}
				#wrapper {
					width: 100%;
					height: 100%;
				}
				#content {
					width: 600px;
					height: 100%;
					padding: 40px 20px;
					margin: auto;
					background-color: #fff;
					border-left: 1px solid #cccccc;
					border-right: 1px solid #cccccc;
				}
				img#wikialogo {
					width: 50%;
					margin: 0px auto;
					display: block;
				}
				div.links {
					margin-top: 30px;
					font-size: 0.8em;
				}
				div.technical {
					margin-top: 60px;
					font-size: 0.6em;
					color: #777;
				}

			</style>
			<!--[if IE]>
			<script src="http://html5shiv.googlecode.com/svn/trunk/html5.js"></script>
			<![endif]-->
		</head>
		<body>
			<div id="wrapper">
				<div id="content">
					<img src="http://upload.wikimedia.org/wikipedia/commons/1/17/Wikia_Logo.svg" id="wikialogo"/>
					<div class="friendly">
						<h1>We are sorry!</h1>
						<p>This problem is due to poor IP communication between back-end computers, possibly including the Web server at the site you are trying to visit. Before analysing this problem, you should clear your browser cache completely.
If you are surfing the Web and see this problem for all Web sites you try to visit, then either:
</p>
<ul><li> your ISP has a major equipment failure/overload
</li><li> there is something wrong with your internal Internet connection e.g. your firewall is not functioning correctly.
</li></ul>
<p>In the first case, only your ISP can help you. In the second case, you need to fix whatever it is that is preventing you reaching the Internet.</p>
					</div>
					<div class="links">
						For more info and updates check out our <a href="https://twitter.com/Wikia">Twitter Feed</a>.
					</div>
					<div class="technical">
						<h2>Technical explanation for geeks and administrators:</h2>
						<h3>502 Bad Gateaway</h3>
						<p>The server, while acting as a gateway or proxy, received an invalid response from the upstream server it accessed in attempting to fulfill the request.</p>
					</div>
			</div> <!-- #content -->
		</div> <!-- #wrapper -->
	</body>
</html>